module execute_tb();
endmodule
